// Deirmentzoglou Ioannis 10015
// deirmentz@ece.auth.gr

`include "Main_Module.sv" 
`include "Normalization.sv"
`include "Rounding.sv"
`include "Exception_Handling.sv"
`include "multiplication.sv"
`include "fp_mult_top.sv"
`include "Assertions.sv" 

